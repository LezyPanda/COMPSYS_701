
module Nios_System_2A (
	clocks_ref_clk_clk,
	clocks_ref_reset_reset,
	clocks_sdram_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	seg_disp_0_external_connection_export,
	seg_disp_1_external_connection_export,
	seg_disp_2_external_connection_export,
	seg_disp_3_external_connection_export,
	seg_disp_5_external_connection_export,
	seg_disp_4_external_connection_export,
	seg_disp_6_external_connection_export);	

	input		clocks_ref_clk_clk;
	input		clocks_ref_reset_reset;
	output		clocks_sdram_clk_clk;
	output	[12:0]	sdram_wire_addr;
	output	[1:0]	sdram_wire_ba;
	output		sdram_wire_cas_n;
	output		sdram_wire_cke;
	output		sdram_wire_cs_n;
	inout	[15:0]	sdram_wire_dq;
	output	[1:0]	sdram_wire_dqm;
	output		sdram_wire_ras_n;
	output		sdram_wire_we_n;
	output	[6:0]	seg_disp_0_external_connection_export;
	output	[6:0]	seg_disp_1_external_connection_export;
	output	[6:0]	seg_disp_2_external_connection_export;
	output	[6:0]	seg_disp_3_external_connection_export;
	output	[6:0]	seg_disp_5_external_connection_export;
	output	[6:0]	seg_disp_4_external_connection_export;
	output	[6:0]	seg_disp_6_external_connection_export;
endmodule
