library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package signal_rom_pkg is
  constant ROM_DEPTH : integer := 1601;
  type rom_t is array (1 to ROM_DEPTH) of std_logic_vector(7 downto 0);
  constant SIGNAL_ROM : rom_t := (
    x"FB",
    x"FF",
    x"F7",
    x"FE",
    x"FC",
    x"F8",
    x"F8",
    x"F8",
    x"FC",
    x"F7",
    x"EA",
    x"EF",
    x"E5",
    x"DE",
    x"DA",
    x"D2",
    x"CB",
    x"C8",
    x"C0",
    x"B9",
    x"B1",
    x"A6",
    x"A2",
    x"9D",
    x"94",
    x"8F",
    x"88",
    x"7F",
    x"7B",
    x"73",
    x"72",
    x"69",
    x"65",
    x"61",
    x"59",
    x"5F",
    x"5A",
    x"55",
    x"56",
    x"4E",
    x"4F",
    x"4C",
    x"4C",
    x"4A",
    x"46",
    x"45",
    x"43",
    x"43",
    x"43",
    x"41",
    x"3B",
    x"3B",
    x"37",
    x"35",
    x"36",
    x"37",
    x"31",
    x"32",
    x"2F",
    x"30",
    x"2A",
    x"2B",
    x"2B",
    x"2B",
    x"2B",
    x"27",
    x"23",
    x"24",
    x"22",
    x"29",
    x"22",
    x"25",
    x"22",
    x"24",
    x"20",
    x"1F",
    x"1E",
    x"22",
    x"20",
    x"20",
    x"23",
    x"20",
    x"20",
    x"22",
    x"1D",
    x"1F",
    x"1F",
    x"1D",
    x"1D",
    x"1A",
    x"1A",
    x"1D",
    x"1E",
    x"22",
    x"1B",
    x"1D",
    x"1D",
    x"19",
    x"1D",
    x"1B",
    x"21",
    x"1E",
    x"20",
    x"20",
    x"22",
    x"21",
    x"24",
    x"26",
    x"28",
    x"25",
    x"22",
    x"25",
    x"2A",
    x"25",
    x"2A",
    x"28",
    x"2B",
    x"24",
    x"28",
    x"26",
    x"2E",
    x"2A",
    x"2C",
    x"27",
    x"28",
    x"29",
    x"2C",
    x"29",
    x"2C",
    x"26",
    x"2A",
    x"2A",
    x"29",
    x"2D",
    x"2D",
    x"2D",
    x"2B",
    x"30",
    x"2E",
    x"2D",
    x"2D",
    x"2C",
    x"28",
    x"2A",
    x"28",
    x"26",
    x"24",
    x"23",
    x"1E",
    x"22",
    x"1E",
    x"1A",
    x"17",
    x"13",
    x"14",
    x"0F",
    x"0B",
    x"0D",
    x"07",
    x"05",
    x"04",
    x"01",
    x"00",
    x"07",
    x"06",
    x"04",
    x"03",
    x"05",
    x"0A",
    x"0F",
    x"0E",
    x"11",
    x"18",
    x"21",
    x"27",
    x"2D",
    x"33",
    x"3A",
    x"40",
    x"4A",
    x"4C",
    x"57",
    x"5C",
    x"64",
    x"6C",
    x"74",
    x"76",
    x"81",
    x"85",
    x"89",
    x"8E",
    x"93",
    x"97",
    x"9B",
    x"9F",
    x"A4",
    x"A8",
    x"A9",
    x"AA",
    x"AE",
    x"B0",
    x"AF",
    x"B5",
    x"B6",
    x"B7",
    x"BA",
    x"BB",
    x"BA",
    x"BE",
    x"BF",
    x"C0",
    x"C7",
    x"C3",
    x"C6",
    x"C7",
    x"C8",
    x"CB",
    x"CD",
    x"D2",
    x"D0",
    x"D0",
    x"D7",
    x"D7",
    x"D5",
    x"D4",
    x"D7",
    x"D8",
    x"DA",
    x"D9",
    x"DB",
    x"DC",
    x"D9",
    x"DA",
    x"DA",
    x"DB",
    x"DC",
    x"DD",
    x"D7",
    x"DD",
    x"E0",
    x"DC",
    x"E1",
    x"E0",
    x"DF",
    x"E0",
    x"DD",
    x"E0",
    x"E4",
    x"E1",
    x"E2",
    x"E0",
    x"E2",
    x"E2",
    x"E3",
    x"E1",
    x"E1",
    x"E5",
    x"DC",
    x"E5",
    x"E1",
    x"E1",
    x"DB",
    x"DD",
    x"DD",
    x"DD",
    x"D8",
    x"DC",
    x"D8",
    x"DA",
    x"DA",
    x"D9",
    x"DA",
    x"D9",
    x"D6",
    x"D7",
    x"D4",
    x"D4",
    x"D8",
    x"D6",
    x"D6",
    x"D8",
    x"D7",
    x"D6",
    x"D8",
    x"D7",
    x"D6",
    x"D3",
    x"D3",
    x"D7",
    x"D0",
    x"D3",
    x"CF",
    x"D5",
    x"D4",
    x"D2",
    x"D1",
    x"CC",
    x"D2",
    x"CC",
    x"CC",
    x"D1",
    x"D0",
    x"D3",
    x"D5",
    x"D7",
    x"D5",
    x"D9",
    x"DA",
    x"DE",
    x"E0",
    x"E3",
    x"E4",
    x"E6",
    x"EC",
    x"E8",
    x"EE",
    x"EF",
    x"F3",
    x"F8",
    x"FA",
    x"F8",
    x"FA",
    x"FC",
    x"FB",
    x"FC",
    x"FB",
    x"F7",
    x"F7",
    x"F0",
    x"F3",
    x"EC",
    x"E6",
    x"E3",
    x"DB",
    x"D8",
    x"D1",
    x"D0",
    x"C7",
    x"B8",
    x"B7",
    x"AC",
    x"A8",
    x"A1",
    x"9B",
    x"93",
    x"90",
    x"85",
    x"81",
    x"7C",
    x"75",
    x"72",
    x"6C",
    x"65",
    x"5F",
    x"63",
    x"5B",
    x"59",
    x"57",
    x"54",
    x"4F",
    x"4E",
    x"4D",
    x"4E",
    x"47",
    x"49",
    x"46",
    x"43",
    x"40",
    x"40",
    x"3E",
    x"3A",
    x"3B",
    x"38",
    x"37",
    x"36",
    x"32",
    x"32",
    x"31",
    x"2B",
    x"30",
    x"31",
    x"2D",
    x"29",
    x"2A",
    x"25",
    x"2B",
    x"28",
    x"27",
    x"23",
    x"25",
    x"22",
    x"22",
    x"22",
    x"20",
    x"20",
    x"21",
    x"1E",
    x"22",
    x"20",
    x"22",
    x"21",
    x"21",
    x"1C",
    x"1D",
    x"1E",
    x"1E",
    x"20",
    x"1D",
    x"20",
    x"1E",
    x"1F",
    x"1D",
    x"1B",
    x"19",
    x"1D",
    x"1E",
    x"1C",
    x"1C",
    x"1D",
    x"1C",
    x"1E",
    x"1F",
    x"20",
    x"21",
    x"23",
    x"23",
    x"27",
    x"25",
    x"28",
    x"24",
    x"27",
    x"26",
    x"28",
    x"28",
    x"23",
    x"25",
    x"25",
    x"29",
    x"2B",
    x"28",
    x"2A",
    x"2A",
    x"27",
    x"2A",
    x"27",
    x"2C",
    x"29",
    x"2D",
    x"29",
    x"2C",
    x"2B",
    x"27",
    x"2A",
    x"2E",
    x"2D",
    x"2B",
    x"2C",
    x"2E",
    x"2B",
    x"2F",
    x"2C",
    x"30",
    x"2A",
    x"2B",
    x"26",
    x"27",
    x"25",
    x"25",
    x"24",
    x"20",
    x"1C",
    x"1C",
    x"19",
    x"15",
    x"13",
    x"10",
    x"0A",
    x"0C",
    x"06",
    x"05",
    x"05",
    x"03",
    x"02",
    x"04",
    x"05",
    x"03",
    x"06",
    x"07",
    x"0A",
    x"0E",
    x"10",
    x"16",
    x"1C",
    x"20",
    x"2A",
    x"2B",
    x"31",
    x"36",
    x"43",
    x"4A",
    x"4F",
    x"58",
    x"5E",
    x"65",
    x"6B",
    x"73",
    x"78",
    x"84",
    x"81",
    x"85",
    x"8C",
    x"91",
    x"96",
    x"9B",
    x"9E",
    x"A3",
    x"A6",
    x"AA",
    x"AE",
    x"B0",
    x"AD",
    x"AD",
    x"B5",
    x"B1",
    x"B7",
    x"B9",
    x"BF",
    x"BC",
    x"BD",
    x"C0",
    x"C2",
    x"C3",
    x"C4",
    x"C4",
    x"C9",
    x"C7",
    x"CA",
    x"D0",
    x"CE",
    x"D0",
    x"D4",
    x"D3",
    x"D7",
    x"D5",
    x"D9",
    x"D9",
    x"D8",
    x"D7",
    x"D8",
    x"DA",
    x"DA",
    x"DA",
    x"DE",
    x"DB",
    x"DF",
    x"DB",
    x"DF",
    x"DC",
    x"DE",
    x"E0",
    x"DD",
    x"DE",
    x"E3",
    x"E1",
    x"DF",
    x"E2",
    x"E0",
    x"E2",
    x"E4",
    x"DE",
    x"E4",
    x"E5",
    x"E2",
    x"E6",
    x"E2",
    x"DF",
    x"DD",
    x"E0",
    x"E2",
    x"E1",
    x"E0",
    x"DD",
    x"DE",
    x"DA",
    x"DB",
    x"DA",
    x"DC",
    x"DA",
    x"D7",
    x"D9",
    x"D7",
    x"D6",
    x"D9",
    x"D7",
    x"D8",
    x"D8",
    x"D7",
    x"D7",
    x"D7",
    x"D8",
    x"D7",
    x"D9",
    x"D6",
    x"D5",
    x"D9",
    x"D4",
    x"D5",
    x"D6",
    x"D4",
    x"D7",
    x"D5",
    x"D4",
    x"D1",
    x"D3",
    x"CF",
    x"D2",
    x"D3",
    x"D1",
    x"D3",
    x"D5",
    x"D3",
    x"D2",
    x"D4",
    x"D4",
    x"D2",
    x"D5",
    x"DB",
    x"DA",
    x"DD",
    x"DD",
    x"E1",
    x"E5",
    x"E4",
    x"EA",
    x"EC",
    x"ED",
    x"F2",
    x"F0",
    x"F2",
    x"F6",
    x"F8",
    x"F9",
    x"F8",
    x"FD",
    x"F8",
    x"FB",
    x"FB",
    x"F7",
    x"F4",
    x"F0",
    x"EA",
    x"E8",
    x"E6",
    x"E2",
    x"D7",
    x"CF",
    x"CC",
    x"C5",
    x"BD",
    x"B4",
    x"B3",
    x"A3",
    x"A0",
    x"97",
    x"92",
    x"8D",
    x"86",
    x"7F",
    x"7C",
    x"76",
    x"71",
    x"6A",
    x"69",
    x"64",
    x"64",
    x"5E",
    x"5B",
    x"56",
    x"51",
    x"50",
    x"4D",
    x"4C",
    x"4C",
    x"48",
    x"45",
    x"45",
    x"43",
    x"43",
    x"3E",
    x"3F",
    x"3D",
    x"3E",
    x"39",
    x"37",
    x"33",
    x"31",
    x"33",
    x"30",
    x"30",
    x"2C",
    x"30",
    x"2B",
    x"2C",
    x"28",
    x"27",
    x"28",
    x"27",
    x"23",
    x"21",
    x"22",
    x"21",
    x"23",
    x"22",
    x"22",
    x"1F",
    x"23",
    x"22",
    x"21",
    x"23",
    x"1F",
    x"21",
    x"20",
    x"20",
    x"1D",
    x"1F",
    x"1D",
    x"1C",
    x"1B",
    x"1F",
    x"1B",
    x"1C",
    x"1A",
    x"1C",
    x"16",
    x"1A",
    x"1A",
    x"1B",
    x"1D",
    x"1D",
    x"22",
    x"1E",
    x"1F",
    x"1D",
    x"20",
    x"1F",
    x"23",
    x"25",
    x"25",
    x"23",
    x"22",
    x"29",
    x"2B",
    x"27",
    x"25",
    x"2A",
    x"27",
    x"27",
    x"2A",
    x"25",
    x"24",
    x"29",
    x"29",
    x"29",
    x"2A",
    x"2B",
    x"2B",
    x"28",
    x"2B",
    x"2A",
    x"29",
    x"28",
    x"2D",
    x"2B",
    x"2C",
    x"2B",
    x"2A",
    x"2E",
    x"2D",
    x"30",
    x"2F",
    x"2F",
    x"2B",
    x"2A",
    x"28",
    x"2B",
    x"2E",
    x"28",
    x"23",
    x"24",
    x"1D",
    x"1A",
    x"1C",
    x"16",
    x"15",
    x"15",
    x"10",
    x"0E",
    x"07",
    x"09",
    x"0A",
    x"05",
    x"00",
    x"02",
    x"01",
    x"03",
    x"04",
    x"06",
    x"07",
    x"09",
    x"0C",
    x"13",
    x"12",
    x"1A",
    x"21",
    x"25",
    x"2D",
    x"33",
    x"38",
    x"41",
    x"47",
    x"4E",
    x"55",
    x"5D",
    x"61",
    x"6A",
    x"71",
    x"76",
    x"7F",
    x"82",
    x"8A",
    x"90",
    x"93",
    x"98",
    x"9D",
    x"9F",
    x"A3",
    x"A3",
    x"AA",
    x"A9",
    x"A9",
    x"B2",
    x"B1",
    x"B4",
    x"B4",
    x"B5",
    x"B2",
    x"BC",
    x"BC",
    x"BE",
    x"C0",
    x"BF",
    x"C2",
    x"C7",
    x"C8",
    x"C6",
    x"C6",
    x"CB",
    x"CE",
    x"D1",
    x"D1",
    x"D0",
    x"D4",
    x"D2",
    x"D4",
    x"D5",
    x"D5",
    x"D8",
    x"D7",
    x"D9",
    x"D9",
    x"DA",
    x"DA",
    x"DE",
    x"DD",
    x"DC",
    x"DA",
    x"DA",
    x"D9",
    x"E3",
    x"E0",
    x"DF",
    x"DD",
    x"DD",
    x"E1",
    x"E3",
    x"DD",
    x"E0",
    x"E1",
    x"DD",
    x"E3",
    x"E1",
    x"E6",
    x"E1",
    x"E3",
    x"DF",
    x"E0",
    x"DF",
    x"E2",
    x"E3",
    x"DF",
    x"E0",
    x"DE",
    x"DE",
    x"E0",
    x"DD",
    x"DA",
    x"D9",
    x"DA",
    x"D9",
    x"D7",
    x"D9",
    x"DA",
    x"D7",
    x"D7",
    x"D2",
    x"D5",
    x"D3",
    x"D5",
    x"D7",
    x"D9",
    x"D9",
    x"D5",
    x"D5",
    x"D7",
    x"D6",
    x"D7",
    x"D6",
    x"D1",
    x"D5",
    x"D4",
    x"D2",
    x"D1",
    x"D5",
    x"D0",
    x"CF",
    x"D2",
    x"D5",
    x"D1",
    x"D1",
    x"CF",
    x"D5",
    x"D2",
    x"D4",
    x"D2",
    x"D7",
    x"D7",
    x"D6",
    x"DA",
    x"DB",
    x"DF",
    x"E1",
    x"E4",
    x"E5",
    x"E9",
    x"EE",
    x"F3",
    x"EF",
    x"F9",
    x"FA",
    x"F9",
    x"F9",
    x"FA",
    x"FD",
    x"FB",
    x"FB",
    x"FC",
    x"FA",
    x"F9",
    x"F5",
    x"F0",
    x"EC",
    x"EA",
    x"E2",
    x"E1",
    x"DA",
    x"D3",
    x"CB",
    x"C5",
    x"C5",
    x"B6",
    x"AC",
    x"AC",
    x"A2",
    x"99",
    x"98",
    x"8E",
    x"87",
    x"7F",
    x"78",
    x"71",
    x"6F",
    x"69",
    x"68",
    x"62",
    x"63",
    x"5F",
    x"59",
    x"56",
    x"56",
    x"4F",
    x"50",
    x"4C",
    x"4A",
    x"48",
    x"48",
    x"44",
    x"42",
    x"43",
    x"3F",
    x"3F",
    x"3C",
    x"3C",
    x"34",
    x"39",
    x"3A",
    x"36",
    x"34",
    x"30",
    x"30",
    x"2E",
    x"2C",
    x"29",
    x"29",
    x"28",
    x"27",
    x"28",
    x"2B",
    x"22",
    x"25",
    x"21",
    x"26",
    x"26",
    x"1F",
    x"26",
    x"20",
    x"22",
    x"24",
    x"21",
    x"25",
    x"26",
    x"20",
    x"1C",
    x"1E",
    x"1D",
    x"1D",
    x"1C",
    x"1E",
    x"22",
    x"1C",
    x"1C",
    x"1F",
    x"1F",
    x"1D",
    x"1E",
    x"1E",
    x"1C",
    x"1E",
    x"1D",
    x"1C",
    x"20",
    x"1F",
    x"1F",
    x"21",
    x"23",
    x"23",
    x"23",
    x"24",
    x"24",
    x"23",
    x"27",
    x"29",
    x"25",
    x"2B",
    x"27",
    x"27",
    x"26",
    x"26",
    x"26",
    x"29",
    x"2C",
    x"2A",
    x"2A",
    x"2B",
    x"24",
    x"29",
    x"2A",
    x"2B",
    x"27",
    x"28",
    x"2C",
    x"2B",
    x"2C",
    x"2A",
    x"29",
    x"2E",
    x"2F",
    x"31",
    x"2A",
    x"2B",
    x"2A",
    x"2D",
    x"2B",
    x"2E",
    x"28",
    x"26",
    x"28",
    x"29",
    x"23",
    x"1F",
    x"1F",
    x"1A",
    x"1A",
    x"19",
    x"15",
    x"0E",
    x"0E",
    x"0C",
    x"0E",
    x"0A",
    x"06",
    x"07",
    x"01",
    x"02",
    x"05",
    x"06",
    x"05",
    x"06",
    x"06",
    x"0C",
    x"0C",
    x"12",
    x"16",
    x"1D",
    x"1F",
    x"27",
    x"2E",
    x"31",
    x"3A",
    x"44",
    x"48",
    x"4E",
    x"57",
    x"5D",
    x"65",
    x"6B",
    x"72",
    x"79",
    x"81",
    x"85",
    x"8D",
    x"8A",
    x"92",
    x"98",
    x"9A",
    x"9C",
    x"A4",
    x"A7",
    x"A9",
    x"AB",
    x"AB",
    x"AE",
    x"B1",
    x"B2",
    x"B6",
    x"BC",
    x"B8",
    x"BC",
    x"BA",
    x"C1",
    x"BE",
    x"C2",
    x"C2",
    x"C6",
    x"C7",
    x"C8",
    x"D0",
    x"CB",
    x"CD",
    x"D5",
    x"CE",
    x"D3",
    x"D1",
    x"D7",
    x"D6",
    x"D8",
    x"D7",
    x"D9",
    x"DC",
    x"D5",
    x"D7",
    x"DC",
    x"DA",
    x"DB",
    x"D9",
    x"DA",
    x"DC",
    x"DB",
    x"DB",
    x"DD",
    x"DC",
    x"E1",
    x"DD",
    x"E3",
    x"DF",
    x"DD",
    x"DF",
    x"E3",
    x"E3",
    x"E2",
    x"E2",
    x"E3",
    x"DF",
    x"E1",
    x"DE",
    x"E1",
    x"E4",
    x"E3",
    x"E6",
    x"E1",
    x"DC",
    x"E3",
    x"E1",
    x"DD",
    x"DE",
    x"DE",
    x"DC",
    x"DC",
    x"DA",
    x"D9",
    x"D9",
    x"D7",
    x"DB",
    x"D7",
    x"D8",
    x"D5",
    x"D4",
    x"D6",
    x"D6",
    x"D8",
    x"D7",
    x"D7",
    x"D3",
    x"D4",
    x"D6",
    x"D5",
    x"D8",
    x"D8",
    x"D3",
    x"D6",
    x"D7",
    x"D4",
    x"D6",
    x"D5",
    x"D2",
    x"D3",
    x"D2",
    x"D0",
    x"D2",
    x"D1",
    x"D0",
    x"D5",
    x"D2",
    x"D8",
    x"D3",
    x"D6",
    x"DA",
    x"DE",
    x"DB",
    x"DB",
    x"E0",
    x"DE",
    x"E3",
    x"E7",
    x"ED",
    x"EF",
    x"EF",
    x"F4",
    x"F4",
    x"F8",
    x"FC",
    x"FA",
    x"FA",
    x"FB",
    x"FD",
    x"FE",
    x"FF",
    x"F9",
    x"F7",
    x"F3",
    x"F4",
    x"ED",
    x"E8",
    x"E8",
    x"E0",
    x"DA",
    x"D0",
    x"CC",
    x"C6",
    x"BB",
    x"B6",
    x"AE",
    x"A9",
    x"9F",
    x"9C",
    x"97",
    x"8C",
    x"86",
    x"81",
    x"7D",
    x"76",
    x"71",
    x"6A",
    x"66",
    x"64",
    x"63",
    x"5D",
    x"56",
    x"57",
    x"53",
    x"51",
    x"4F",
    x"4B",
    x"4A",
    x"48",
    x"47",
    x"46",
    x"44",
    x"42",
    x"40",
    x"3F",
    x"3E",
    x"3E",
    x"3B",
    x"37",
    x"37",
    x"34",
    x"2F",
    x"2C",
    x"2C",
    x"2D",
    x"2B",
    x"2A",
    x"2A",
    x"27",
    x"26",
    x"28",
    x"27",
    x"2A",
    x"25",
    x"24",
    x"22",
    x"23",
    x"23",
    x"1F",
    x"21",
    x"23",
    x"20",
    x"22",
    x"23",
    x"23",
    x"22",
    x"1B",
    x"1E",
    x"21",
    x"1F",
    x"1E",
    x"1F",
    x"20",
    x"1D",
    x"1B",
    x"1C",
    x"1C",
    x"1E",
    x"1D",
    x"1E",
    x"1D",
    x"1C",
    x"1D",
    x"1E",
    x"1B",
    x"1F",
    x"21",
    x"20",
    x"24",
    x"23",
    x"22",
    x"23",
    x"23",
    x"25",
    x"27",
    x"25",
    x"27",
    x"2A",
    x"29",
    x"29",
    x"26",
    x"27",
    x"29",
    x"28",
    x"25",
    x"25",
    x"2B",
    x"27",
    x"2D",
    x"24",
    x"2A",
    x"29",
    x"28",
    x"2B",
    x"29",
    x"2D",
    x"2B",
    x"28",
    x"27",
    x"2C",
    x"2F",
    x"2E",
    x"2E",
    x"2F",
    x"2A",
    x"30",
    x"2B",
    x"2C",
    x"2A",
    x"2A",
    x"24",
    x"29",
    x"25",
    x"26",
    x"23",
    x"1D",
    x"18",
    x"14",
    x"15",
    x"12",
    x"11",
    x"0B",
    x"0C",
    x"08",
    x"04",
    x"06",
    x"04",
    x"02",
    x"06",
    x"04",
    x"03",
    x"06",
    x"07",
    x"0A",
    x"0E",
    x"10",
    x"14",
    x"1B",
    x"24",
    x"25",
    x"2A",
    x"32",
    x"39",
    x"40",
    x"49",
    x"4F",
    x"55",
    x"5C",
    x"62",
    x"69",
    x"6F",
    x"77",
    x"7C",
    x"82",
    x"89",
    x"8C",
    x"93",
    x"98",
    x"99",
    x"A1",
    x"9F",
    x"A5",
    x"A5",
    x"AA",
    x"AA",
    x"AE",
    x"B0",
    x"B1",
    x"B1",
    x"B8",
    x"BD",
    x"BF",
    x"BB",
    x"BE",
    x"BF",
    x"C2",
    x"C1",
    x"C1",
    x"C7",
    x"C6",
    x"C6",
    x"D1",
    x"CD",
    x"D0",
    x"D3",
    x"CE",
    x"D4",
    x"D6",
    x"D6",
    x"D7",
    x"D6",
    x"DA",
    x"D7",
    x"D8",
    x"DC",
    x"DE",
    x"DA",
    x"DB",
    x"DD",
    x"DE",
    x"DF",
    x"DD",
    x"DC",
    x"DF",
    x"DE",
    x"E1",
    x"DC",
    x"DF",
    x"E2",
    x"DF",
    x"DF",
    x"DF",
    x"E0",
    x"E1",
    x"E2",
    x"E0",
    x"E2",
    x"E1",
    x"E1",
    x"E0",
    x"E1",
    x"E9",
    x"E8",
    x"E3",
    x"E2",
    x"DD",
    x"DD",
    x"DD",
    x"DE",
    x"DD",
    x"DC",
    x"DA",
    x"D8",
    x"DA",
    x"DB",
    x"D9",
    x"D8",
    x"D9",
    x"D8",
    x"D3",
    x"D6",
    x"D5",
    x"D2",
    x"D3",
    x"D5",
    x"D7",
    x"D5",
    x"D6",
    x"D4",
    x"D1",
    x"D5",
    x"D3",
    x"D7",
    x"D8",
    x"D3",
    x"D6",
    x"D5",
    x"D0",
    x"D2",
    x"D2",
    x"D2",
    x"D2",
    x"D2",
    x"D2",
    x"D0",
    x"D2",
    x"CD",
    x"D0",
    x"D6",
    x"D3",
    x"D7",
    x"DB",
    x"D8",
    x"DA",
    x"DE",
    x"E2",
    x"E3",
    x"E5",
    x"E6",
    x"EC",
    x"EF",
    x"F1",
    x"F4",
    x"F4",
    x"FA",
    x"F5"
  );
end package signal_rom_pkg;
